* /home/pavan.gutti2/Desktop/pavang_cla_adder/pavang_cla_adder.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sat 05 Mar 2022 03:51:20 PM UTC

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U18  Net-_U12-Pad10_ Net-_U12-Pad11_ Net-_U12-Pad12_ Net-_U12-Pad13_ Net-_U12-Pad14_ o0 o1 o2 o3 o4 dac_bridge_5		
U12  Net-_U10-Pad5_ Net-_U10-Pad6_ Net-_U10-Pad7_ Net-_U10-Pad8_ Net-_U11-Pad6_ Net-_U11-Pad7_ Net-_U11-Pad8_ Net-_U11-Pad9_ Net-_U11-Pad10_ Net-_U12-Pad10_ Net-_U12-Pad11_ Net-_U12-Pad12_ Net-_U12-Pad13_ Net-_U12-Pad14_ pavan_cla_adder		
U10  i0 i1 i2 i3 Net-_U10-Pad5_ Net-_U10-Pad6_ Net-_U10-Pad7_ Net-_U10-Pad8_ adc_bridge_4		
U11  i4 i5 i6 i7 i8 Net-_U11-Pad6_ Net-_U11-Pad7_ Net-_U11-Pad8_ Net-_U11-Pad9_ Net-_U11-Pad10_ adc_bridge_5		
v0  i0 GND pulse		
v1  i1 GND pulse		
v2  i2 GND pulse		
v3  i3 GND pulse		
v7  i7 GND pulse		
v6  i6 GND pulse		
v5  i5 GND pulse		
v4  i4 GND pulse		
v8  i8 GND pulse		
U5  i4 plot_v1		
U6  i5 plot_v1		
U7  i6 plot_v1		
U9  i8 plot_v1		
U1  i0 plot_v1		
U2  i1 plot_v1		
U3  i2 plot_v1		
U4  i3 plot_v1		
U8  i7 plot_v1		
R1  o0 GND 1k		
R3  o2 GND 1k		
R4  o3 GND 1k		
R5  o4 GND 1k		
R2  o1 GND 1k		
U13  o0 plot_v1		
U14  o1 plot_v1		
U15  o2 plot_v1		
U17  o4 plot_v1		
U16  o3 plot_v1		

.end
